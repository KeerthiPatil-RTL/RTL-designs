module comp4bit_eqn (
    input  [3:0] A, B,
    output G, E, L
);

assign E = (A[3] ~^ B[3]) & 
           (A[2] ~^ B[2]) & 
           (A[1] ~^ B[1]) & 
           (A[0] ~^ B[0]);

assign G = (A[3] & ~B[3]) |
           (A[2] & ~B[2] & (A[3] ~^ B[3])) |
           (A[1] & ~B[1] & (A[3] ~^ B[3]) & (A[2] ~^ B[2])) |
           (A[0] & ~B[0] & (A[3] ~^ B[3]) & (A[2] ~^ B[2]) & (A[1] ~^ B[1]));

assign L = (~A[3] & B[3]) |
           (~A[2] & B[2] & (A[3] ~^ B[3])) |
           (~A[1] & B[1] & (A[3] ~^ B[3]) & (A[2] ~^ B[2])) |
           (~A[0] & B[0] & (A[3] ~^ B[3]) & (A[2] ~^ B[2]) & (A[1] ~^ B[1]));

endmodule

